module DataMemory(clk, Address, WriteData, MemWrite, MemRead, ReadData);

reg [7:0] Memory [0:1023];



endmodule
