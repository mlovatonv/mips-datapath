module DataMemory(clk, Address, WriteData, ReadData);
